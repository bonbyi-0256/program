module selector8_tb;
  reg [2:0] s;
  reg [0:7] a;
  wire x;

  selector8 selector8_0(.s(s),.a(a),.x(x));

  initial begin
  $dumpvars;
  s=7;
  a=8'b00000000;#100
  a=8'b00000001;#100
  a=8'b00000010;#100
  a=8'b00000011;#100
  a=8'b00000100;#100
  a=8'b00000111;#100
  a=8'b00001000;#100
  a=8'b00001111;#100
  a=8'b00010000;#100
  a=8'b00011111;#100
  a=8'b00100000;#100
  a=8'b00111111;#100
  a=8'b01000000;#100
  a=8'b01111111;#100
  a=8'b10000000;#100
  a=8'b11111111;#100
  $finish;
  end

endmodule